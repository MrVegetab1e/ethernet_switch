`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/06/29 15:01:48
// Design Name: 
// Module Name: hash_tte_bucket
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
//====================================================================
//entry structure:
//[15:0]:portmap
//[63:16]:dst mac
//[111:64]:src mac
//[119]:item valid
//=====================================================================
module hash_tte_bucket(
input               clk,
input               rstn,
//port se signals.
input       [47:0]  se_dmac,
input       [47:0]  se_smac, ///用于流表匹配时的源mac地址
input       [11:0]  se_hash,        
input               se_req,
output  reg         se_ack,
output  reg         se_nak,
output  reg [15:0]  se_result,
input               hash_clear, ///清空ram
input               hash_update, ////更新ram
input       [11:0]  hash,
input       [119:0] flow,
output  reg         reg_rst    ////插入流表成功后返回1
);
//======================================
//              main state.
//======================================

reg     [2:0]   state;
reg             clear_op;
// reg             hit;
reg     [1:0]   hit_0, hit_1;
wire            item_valid;
//======================================
//              one cycle for state1.
//======================================
reg     [ 1:0]  count;

reg     [47:0]  hit_dmac;
reg     [47:0]  hit_smac;

// reg             init;
reg                 ram_wr;
reg     [11:0]      ram_addr;     //input  [11 : 0] addra
reg     [119:0]     ram_din;      //input  [119 : 0] dina
wire    [119:0]     ram_dout;     //output [119 : 0] douta
// reg     [119:0]     ram_dout_reg; //output [119 : 0] douta


parameter   HASH0 = 12'b0110_1000_1110;
parameter   DEST_MAC0 =48'h60beb403060e;
parameter   SOURCE_MAC0 = 48'h60beb403644d;
parameter   HASH_PORT0 = 16'b0010;
parameter   HASH_VALID0 = 8'b10000000;

parameter   HASH1 = 12'b0111_0100_1101;
parameter   DEST_MAC1 =48'h60beb403644d;
parameter   SOURCE_MAC1 = 48'h60beb403060e;
parameter   HASH_PORT1 = 16'b0100;
parameter   HASH_VALID1 = 8'b10000000;

always @(posedge clk or negedge rstn)
    if(!rstn) begin
        state <=#2 0;
        // init <=#2 0;
        clear_op<=#2 1;
        ram_wr<=#2 0;
        ram_addr<=#2 0; 
        // ram_din<=#2 0;     
        se_ack<=#2 0;
        se_nak<=#2 0;
        // se_result<=#2 0;
        // hit_dmac<=#2 0;
        // hit_smac<=#2 0;
        hit_0<=#2 0;
        hit_1<=#2 0;
        count<=#2 0;
        reg_rst<=#2 0;
        end
    else begin
        // ram_dout_reg<=#2 ram_dout;
        ram_wr<=#2 0;
        se_ack<=#2 0;
        se_nak<=#2 0;
        // reg_rst<=#2 0;
        // ram_din<=#2 flow; 
        case(state)
            0:begin
                if(hash_clear | clear_op)begin
                    ram_addr<=#2 0;   
                    ram_wr<=#2 1;
                    ram_din<=#2 0;
                    state<=#2 6;
                    reg_rst<=#2 1;
                end
                else if(hash_update)begin
                    ram_addr<=#2 hash; 
                    ram_wr<=#2 1;
                    ram_din<=#2 flow; 
                    state<=#2 4;
                    reg_rst<=#2 1;
                end
                else if(se_req) begin
                    ram_addr<=#2 se_hash;
                    hit_dmac   <=#2 se_dmac;
                    hit_smac   <=#2 se_smac;
                    count     <=#2 0;
                    state   <=#2 1;
                end
                // else if(init) begin
                //     ram_addr<=#2 HASH0;   
                //     ram_wr<=#2 1;
                //     ram_din<=#2 {HASH_VALID0,SOURCE_MAC0,DEST_MAC0,HASH_PORT0};
                //     state<=#2 7; 
                // end
            end
            1:begin
                // count <=#2 1;
                // if(count) state<=#2 2;
                count <=#2 {count, 1'b1};
                if(count[1]) state<=#2 2;
            end
            2:begin
                hit_0<={hit_dmac[0+:24]==ram_dout[16+:24], hit_dmac[24+:24]==ram_dout[40+:24]};
                hit_1<={hit_smac[0+:24]==ram_dout[64+:24], hit_smac[24+:24]==ram_dout[88+:24]};
                se_result<=#2 ram_dout[15:0];
                state<=#2 3;
            end
            3:begin
                // if(hit)begin
                if((hit_0 == 2'b11) && (hit_1 == 2'b11) && item_valid) begin
                    se_nak<=#2 0;
                    se_ack<=#2 1;
                    // se_result<=#2 ram_dout_reg[15:0];
                end
                else begin
                    se_ack<=#2 0;
                    se_nak<=#2 1;
                end
                state<=#2 5;
            end
            4:begin
                reg_rst<=#2 0;
                state<=#2 0;
            end
            5:begin
                state<=#2 0;
            end
            6:begin
                if(ram_addr<12'hfff) begin
                    ram_addr<=#2 ram_addr+1;
                    ram_wr<=#2 1;
                end
                else begin
                    ram_addr<=#2 0;
                    ram_wr<=#2 0;
                    clear_op<=#2 0;
                    reg_rst<=#2 0;
                    state<=#2 0;
                end
            end
            // 7:begin
            //     ram_addr<=#2 HASH1;   
            //     ram_wr<=#2 1;
            //     ram_din<=#2 {HASH_VALID1,SOURCE_MAC1,DEST_MAC1,HASH_PORT1};
            //     init <=#2 0;
            //     state<=#2 0;
            // end
        endcase
    end 

// always @(*)begin
//     hit=(hit_dmac==ram_dout_reg[63:16])&(hit_smac==ram_dout_reg[111:64])&item_valid;                   
//     end
//assign item_valid=ram_dout_reg[119];
assign item_valid = ram_dout[119];

sram_reg2_w120_d4k u_sram_0 (
  .clka(clk),           // input clka
  .wea(ram_wr),       // input  [0 : 0] wea
  .addra(ram_addr),   // input  [11 : 0] addra
  .dina(ram_din),     // input  [119 : 0] dina
  .douta(ram_dout)    // output [119 : 0] douta
);

endmodule
